import uvm_pkg::*;
`include "reg_file.sv"
`include "seq_item.sv"
`include "ftm_if.sv"
`include "ftm_if2.sv"
`include "sync_mem.sv"
`include "dut_mem.sv"
`include "sequence.sv"
`include "ftm_seqr.sv"
`include "epwm_reference_sb.sv"
`include "cpwm_reference_sb.sv"
`include "output_compare_reference_sb.sv"
`include "epwm_checker.sv"
`include "cpwm_checker.sv"
`include "output_compare_checker.sv"
`include "calculation_scoreboard.sv"
`include "ftm_driver.sv"
`include "input_monitor.sv"
`include "output_monitor.sv"
`include "ftm_dut.sv"
`include "optcomp_sc.sv"
`include "edgealigned_pwm_sc.sv"
`include "cntralig_sc.sv"
`include "ftm_agent.sv"
`include "ftm_dut_agent.sv"
`include "ftm_env.sv"
`include "ftm_dut_env.sv"
`include "ftm_test.sv"

