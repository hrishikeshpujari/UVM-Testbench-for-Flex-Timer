
interface ftm_if;
 bit CH0;	
 bit CH1;	
 bit CH2;	
 bit CH3;	
 bit CH4;	
 bit CH5;	
 bit CH6;	
 bit CH7;	
 bit [0:31] data;
 bit clk;
 bit wr_en;
 bit rd_en; 
 reg_name_enum reg_name;

 //ftm_sc FTM_SC;
 //ftm_cnt FTM_CNT;
 //ftm_mod FTM_MOD;
 //ftm_csc FTM_CSC;
 //ftm_cnv FTM_CNV;
 //ftm_cntin FTM_CNTIN;
 //ftm_status FTM_STATUS;
 //ftm_mode FTM_MODE;
 //ftm_sync FTM_SYNC;
 //ftm_outinit FTM_OUTINIT;
 //ftm_outmask FTM_OUTMASK;
 //ftm_combine FTM_COMBINE;
 //ftm_deadtime FTM_DEADTIME;
 //ftm_exttrig FTM_EXTTRIG;
 //ftm_pol FTM_POL;
 //ftm_fms FTM_FMS;
 //ftm_filter FTM_FILTER;
 //ftm_qdctrl FTM_QDCTRL;
 //ftm_conf FTM_CONF;
 //ftm_synconf FTM_SYNCONF;
 //ftm_invctrl FTM_INVCTRL;
 //ftm_swoctrl FTM_SWOCTRL;
 //ftm_pwmload FTM_PWMLOAD;

endinterface: ftm_if

